entity attrdecl1 is
end;

architecture behav of attrdecl1 is
  attribute user_attr : string;
begin
end;
