entity stdhide1 is
end;

architecture behav of stdhide1 is
  constant min : natural := 5;
begin
end;
