entity complexstmtlayout4 is
end;

architecture behav of complexstmtlayout4 is
begin
  process
    variable a : boolean;
  begin
    for i in 1 to 5 loop
      null;
    end loop;
  end process;
end behav;
