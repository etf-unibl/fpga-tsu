entity port1 is
  port (data_i : bit;
        data_o : out bit;
        d2_b : inout bit);
end;
