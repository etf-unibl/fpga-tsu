-----------------------------------------------------------------------------
-- This is a correct comment.
-----------------------------------------------------------------------------
-- Also an empty comment
--
