entity generic2 is
  generic (g_bad : natural := 1);
end;
