entity subprgislayout1 is
end;

architecture behav of subprgislayout1 is
begin
  process
    procedure p
    is
      constant c : natural := 5;
    begin
      null;
    end p;
  begin
      null;
  end process;
end behav;
