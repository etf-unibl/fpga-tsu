entity paren4 is
end;

architecture behav of paren4 is
  function f return natural is
  begin
    return 4;
  end f;
begin
end behav;
