entity entitylayout2 is
  generic (
    a : bit := '0';
    b : integer := 2
  );
end;
