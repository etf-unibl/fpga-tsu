entity indent4 is
  type t1 is range 1 to 3;
    type t2 is range 1 to 3;
 subtype t3 is natural range 4 to 5;
end;
