entity entitylayout6 is
  generic (
    a : bit     := '0';
    b : integer := 2
  );
  port (
    i1 :     bit;
    o1 : out bit
  );
end;
