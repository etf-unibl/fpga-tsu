entity reference12 is
  constant c : character := NUL;
end;
  
