library ieee, unisims;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

use work.my_pkg.all;

entity contextclauses4 is
end;
