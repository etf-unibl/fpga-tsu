use std.textio;

entity reference5 is
end;
