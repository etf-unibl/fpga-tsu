library std;
use std.textio.all;

entity contextclauses3 is
end;
