entity complexstmtlayout7 is
end;

architecture behav of complexstmtlayout7 is
begin
  process
    variable a : boolean;
  begin
    while False loop
      null;
    end loop;
  end process;
end behav;
