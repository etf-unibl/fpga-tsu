use std.textio;

entity contextuse1 is
end;
