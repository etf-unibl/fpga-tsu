use std.textio.all;

entity contextclauses1 is
end contextclauses1;
