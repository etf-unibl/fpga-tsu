entity entitylayout3 is
  generic (
    a     : bit;
    b : integer := 2
  );
end;
