entity generic1 is
  generic (g_ONE : natural := 1);
end;
