entity port3 is
  port (v_in : bit);
end;
