entity namedecl1 is
end;

architecture behav of namedecl1 is
  constant Reserved : natural := 5;
begin
end;
