library work;
use work.foo.all;

entity contextclauses2 is
end;
