entity reference17 is
  attribute Attr : natural;
  attribute Attr of reference17 : entity is 5;
end;
