entity signalsname1 is
end;

architecture arch of signalsname1 is
  signal s : bit;
  signal s1_n : bit;
  signal s1_a : bit;
  signal s_p : bit;
begin
end;
