entity operatorspace3 is
  constant c : boolean := 4 >  2;
end;

