library ieee;
use ieee.std_logic_1164.all;

entity porttypes3 is
  port (a : std_ulogic_vector(3 downto 0));
end;
