library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

library unisims;
use unisims.VPKG.all;

library proj_pci;
use proj_pci.pci_defs.all;

use work.my_pkg.all;

entity contextclauses4 is
end;
