entity simpleblock4 is
end;

architecture behav of simpleblock4 is
  signal s : bit;
begin
  b: block
  begin
  end block;
end;
