entity entityitems1 is
  constant c : natural := 5;
end;
