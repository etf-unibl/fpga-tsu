library ieee;

entity dependences3 is
end;


architecture behav of dependences3 is
  use ieee.std_logic_1164.all;
  signal s : std_logic;
begin
  s <= '0';
end;
