entity indent9 is
end;

library ieee;

architecture behav of indent9 is
    use ieee.std_logic_1164.all;
begin
end;
