entity hello is
end;


