use STD.textio;

entity reference6 is
end;
