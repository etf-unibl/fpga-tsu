entity signalsname3 is
end;

architecture arch of signalsname3 is
  signal s_n_a : bit;
begin
end;
