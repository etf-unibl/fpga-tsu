entity attrdecl1 is
end;

architecture behav of attrdecl1 is
  attribute reserved : boolean;
begin
end;
