library ieee;
use ieee.std_logic_1164.all;

entity nospace5 is
end nospace5;
