architecture onemodule2 of onemodule1 is
begin
end;
