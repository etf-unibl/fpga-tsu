--  Incorrect place for generic
entity indent1 is
generic (g : natural);
end indent1;
