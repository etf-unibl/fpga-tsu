entity port2 is
  port (v : out bit);
end;
