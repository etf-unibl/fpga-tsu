entity reference1 is
  generic (g1: natural := 5);
begin
  assert g1 > 2;
end;
