library ieee;
use ieee.std_logic_1164.all;

entity porttypes2 is
  port (a : std_ulogic);
end;
