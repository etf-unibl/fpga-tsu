entity operatorspace1 is
  constant c : integer := 4/ 2;
end;

