entity beginendlayout4 is
end;

architecture behav of beginendlayout4 is
begin
  b : block
    begin
  end block b;
end behav;
