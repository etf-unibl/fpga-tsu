entity beginendlayout3 is
end;

architecture behav of beginendlayout3 is
  begin
end behav;
