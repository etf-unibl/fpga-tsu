entity namedecl2 is
end;

architecture behav of namedecl2 is
  constant ok : natural := 5;
begin
end;
