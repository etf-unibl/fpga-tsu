entity nospace1 is
  constant c :boolean := True;
end nospace1;
