package onemodule4 is
end;

package body onemodule4 is
end;
