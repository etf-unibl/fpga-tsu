-- This file has two lines of exactely 80 characters.
--000000011111111112222222222333333333344444444445555555555666666666677777777778
--345678901234567890123456789012345678901234567890123456789012345678901234567890
