--  Bad character �
entity charset1 is
end;
