library ieee;
use ieee.std_logic_1164.all;

entity reference8 is
  constant c : std_logic := '1';
end;
