entity simpleblock2 is
end;

architecture behav of simpleblock2 is
begin
  b: block
    port (s : bit);
  begin
  end block;
end;
