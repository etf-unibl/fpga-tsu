entity contextuse2 is
  use std.textio;
end;
