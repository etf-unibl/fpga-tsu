entity reference11 is
  constant c : Bit_Vector := "01";
end;
