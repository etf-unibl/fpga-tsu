--This is an incorrect comment (missing space).
entity comment1 is
end;
