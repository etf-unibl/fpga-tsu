entity port4 is
  port (b_o : buffer bit);
end;
