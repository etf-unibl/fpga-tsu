entity beginendlayout8 is
end;

architecture behav of beginendlayout8 is
begin
  process
    procedure p is
      begin
        null;
    end p;
  begin
      null;
  end process;
end behav;
