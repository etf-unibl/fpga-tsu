entity beginendlayout6 is
end;

architecture behav of beginendlayout6 is
begin
  process
    begin
      null;
  end process;
end behav;
