entity beginendlayout1 is
begin
end;
