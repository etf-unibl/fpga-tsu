--  There is a space at the end of this line  
