entity beginendlayout2 is
 begin
end;
