entity ieeepkg1 is
end;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

architecture behav of ieeepkg1 is
  signal s : std_logic;
begin
end;
