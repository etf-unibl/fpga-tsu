entity spaces1 is
  constant c : boolean := 1 >3;
end;
