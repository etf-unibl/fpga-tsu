entity onemodule8 is
end;

architecture behav2 of onemodule8 is
begin
end;

configuration onemodule8_conf of onemodule8 is
  for behav2
  end for;
end;

