entity attrname2 is
end;

architecture behav of attrname2 is
  constant n : string := "hello";
  constant l : natural := n'left;
begin
end;
