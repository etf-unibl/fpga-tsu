package onemodule5 is
end;

package body onemodule4 is
end;
