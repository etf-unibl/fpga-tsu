library Work;

entity reference4 is
end;
