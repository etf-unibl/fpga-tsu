entity endlabel1 is
end;
