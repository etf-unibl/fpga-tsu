entity dependences2 is
end;

library ieee;
use ieee.std_logic_1164.all;

architecture behav of dependences2 is
  signal s : std_logic;
begin
  s <= '0';
end;
