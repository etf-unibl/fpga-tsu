package onemodule7 is
end;

package body onemodule7 is
end;

package onemodule7b is
end;
