entity enum2 is
  type my_enum is (S0, S1, S2, err);
end;
  
