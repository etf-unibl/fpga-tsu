entity complexstmtlayout6 is
end;

architecture behav of complexstmtlayout6 is
begin
  process
    variable a : boolean;
  begin
    for i in 1 to 5
      loop
      null;
    end loop;
  end process;
end behav;
