entity processlabel1 is
end;

architecture behav of processlabel1 is
begin
  tchk: process
  begin
    null;
  end process;
end;
