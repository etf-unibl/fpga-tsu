use std.TEXTIO;

entity reference7 is
end;
