entity entityitems2 is
begin
  process
  begin
    wait;
  end process;
end;
