-- This file is using-- (old) Mac OS newline-- convention. That is \r
