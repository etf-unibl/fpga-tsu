entity signalsname2 is
end;

architecture arch of signalsname2 is
  signal s_o : bit;
begin
end;
