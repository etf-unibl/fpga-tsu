entity beginendlayout7 is
end;

architecture behav of beginendlayout7 is
  function f return natural is
    begin
      return 5;
  end;
begin
  process
  begin
      null;
  end process;
end behav;
