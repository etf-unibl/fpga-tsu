entity reference2 is
  generic (G1: natural := 5);
begin
  assert g1 > 2;
end;
