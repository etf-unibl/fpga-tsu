library ieee;
use ieee.std_logic_1164.all;

entity stdhide2 is
end;

architecture behav of stdhide2 is
  constant std_logic : natural := 5;
begin
end;
