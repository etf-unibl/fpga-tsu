entity onemodule3 is
end;

-- Not ok: unrelated arc

architecture behav2 of onemodule1 is
begin
end;
