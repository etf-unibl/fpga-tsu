library ieee;
use ieee.std_logic_1164.all;

entity dependences1 is
end;

architecture behav of dependences1 is
  signal s : std_logic;
begin
  s <= '0';
end;
