library work;

entity reference3 is
end;
