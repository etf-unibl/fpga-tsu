entity complexstmtlayout8 is
end;

architecture behav of complexstmtlayout8 is
begin
  process
    variable a : boolean;
  begin
    while False
     loop
      null;
    end loop;
  end process;
end behav;
