entity forbiddenid is
  constant l : natural := 1;
end;

