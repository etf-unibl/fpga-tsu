entity processlabel3 is
end;

architecture behav of processlabel3 is
begin
  --  Comment not for the assert.

  process
  begin
    wait;
  end process;
end;
