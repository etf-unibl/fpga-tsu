--- this is a very very very very very very very very very very very very very long line.
