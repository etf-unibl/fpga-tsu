entity onemodule1 is
end;
