entity filename1_err is
end;
