entity operatorspace1 is
  constant c : integer := 1 +3;
end;

