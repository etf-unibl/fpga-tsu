entity entitylayout4 is
  port (
    i1 : in bit := '0';
    o1 : out bit
  );
end;
