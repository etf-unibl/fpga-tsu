entity hello is
end;


