library ieee;
use ieee.std_logic_1164.all;

entity porttypes1 is
  port (a : std_logic;
        b : std_logic_vector(7 downto 0));
end;
