entity indent6 is
end;

architecture behav of indent6 is
  constant b : bit_vector := x"a5";
   attribute attr : natural;
begin
end;
