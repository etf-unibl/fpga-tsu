--  Incorrect place for port
entity indent1 is
port (g : natural);
end indent1;
