entity generic3 is
  generic (BAD : natural := 1);
end;
