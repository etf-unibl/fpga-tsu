entity beginendlayout5 is
end;

architecture behav of beginendlayout5 is
begin
  g : for i in 1 to 2 generate
    begin
  end generate g;
end behav;
