entity enumcharlit1 is
end;

architecture behav of enumcharlit1 is
  type my_enum is (aa, bb, 'c');
begin
end;
