entity dependences3 is
end;

library ieee;

architecture behav of dependences3 is
  signal s : ieee.std_logic_1164.std_logic;
begin
end;
