library ieee;
use ieee.std_logic_1164.all;

entity reference9 is
  constant c : STD_LOGIC := '1';
end;
