entity reference10 is
  constant c : string := "hello";
end;
