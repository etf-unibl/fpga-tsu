package onemodule6 is
end;

package onemodule6b is
end;
