entity nospace5 is
  constant c : character := character' Val(4);
end nospace5;
